// Benchmark "c3540" written by ABC on Thu Aug 22 15:03:06 2019

module c3540 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21;
  wire n73, n74, n76, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n107, n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
    n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
    n140, n141, n142, n143, n144, n145, n146, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n435, n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n553,
    n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
    n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
    n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
    n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
    n724, n725, n726, n727, n728, n729, n730, n731, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
    n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
    n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1004,
    n1005, n1006, n1007, n1008, n1009, n1011, n1012, n1013, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
       n1038, n1039, n1040, n1041, n1042;
  wire po11_prelocked, po12_prelocked, po13_prelocked, po14_prelocked, po15_prelocked, po16_prelocked, po17_prelocked, po18_prelocked, po19_prelocked, po20_prelocked, po21_prelocked;
  wire rest0, rest1, rest2, rest3, rest4, rest5, rest6, rest7, rest8, rest9, rest10, rest11, rest12, rest13, rest14, rest15;
  wire sf_in0_s, sf_in1_s, sf_in2_s, sf_in3_s, sf_in4_s, sf_in5_s, sf_in6_s, sf_in7_s, sf_in8_s, sf_in9_s, sf_in10_s, sf_in11_s, sf_in12_s, sf_in13_s, sf_in14_s;
  wire sf_in0_c, sf_in1_c, sf_in2_c, sf_in3_c, sf_in4_c, sf_in5_c, sf_in6_c, sf_in7_c, sf_in8_c, sf_in9_c, sf_in10_c, sf_in11_c, sf_in12_c, sf_in13_c, sf_in14_c;
  wire rest_in0_s, rest_in1_s, rest_in2_s, rest_in3_s, rest_in4_s, rest_in5_s, rest_in6_s, rest_in7_s, rest_in8_s, rest_in9_s, rest_in10_s, rest_in11_s, rest_in12_s, rest_in13_s, rest_in14_s;
  wire rest_in0_c, rest_in1_c, rest_in2_c, rest_in3_c, rest_in4_c, rest_in5_c, rest_in6_c, rest_in7_c, rest_in8_c, rest_in9_c, rest_in10_c, rest_in11_c, rest_in12_c, rest_in13_c, rest_in14_c;
  wire hd, rest;
  wire sp_in0, sp_in1, sp_in2, sp_in3, sp_in4, sp_in5, sp_in6, sp_in7, sp_in8, sp_in9, sp_in10, sp_in11, sp_in12, sp_in13, sp_in14, sp_in15;
  wire sp_sf_in0, sp_sf_in1, sp_sf_in2, sp_sf_in3, sp_sf_in4, sp_sf_in5, sp_sf_in6, sp_sf_in7, sp_sf_in8, sp_sf_in9, sp_sf_in10, sp_sf_in11, sp_sf_in12, sp_sf_in13, sp_sf_in14, sp_sf_in15;
  

  wire fa_in8_int0, fa_in9_int0, fa_in10_int0, fa_in11_int0;
  wire fa_in8_int1, fa_in9_int1, fa_in10_int1, fa_in11_int1;
  wire fa_in8_int2, fa_in9_int2, fa_in10_int2, fa_in11_int2;
  wire fa_in8_s, fa_in9_s, fa_in10_s, fa_in11_s;
  wire fa_in8_c, fa_in9_c, fa_in10_c, fa_in11_c;
  
  wire fa1_in12_int0, fa1_in13_int0, fa2_in12_int0, fa2_in13_int0;
  wire fa1_in12_int1, fa1_in13_int1, fa2_in12_int1, fa2_in13_int1;
  wire fa1_in12_int2, fa1_in13_int2, fa2_in12_int2, fa2_in13_int2;
  wire fa1_in12_s, fa1_in13_s, fa2_in12_s, fa2_in13_s;
  wire fa1_in12_c, fa1_in13_c, fa2_in12_c, fa2_in13_c;
  
  wire fa1_in14_int0, fa2_in14_int0, fa3_in14_int0;
  wire fa1_in14_int1, fa2_in14_int1, fa3_in14_int1;
  wire fa1_in14_int2, fa2_in14_int2, fa3_in14_int2;
  wire fa1_in14_s, fa2_in14_s, fa3_in14_s;
  wire fa1_in14_c, fa2_in14_c, fa3_in14_c;
  
  wire restfa_in8_int0, restfa_in9_int0, restfa_in10_int0, restfa_in11_int0;
  wire restfa_in8_int1, restfa_in9_int1, restfa_in10_int1, restfa_in11_int1;
  wire restfa_in8_int2, restfa_in9_int2, restfa_in10_int2, restfa_in11_int2;
  wire restfa_in8_s, restfa_in9_s, restfa_in10_s, restfa_in11_s;
  wire restfa_in8_c, restfa_in9_c, restfa_in10_c, restfa_in11_c;
  
  wire restfa1_in12_int0, restfa1_in13_int0, restfa2_in12_int0, restfa2_in13_int0;
  wire restfa1_in12_int1, restfa1_in13_int1, restfa2_in12_int1, restfa2_in13_int1;
  wire restfa1_in12_int2, restfa1_in13_int2, restfa2_in12_int2, restfa2_in13_int2;
  wire restfa1_in12_s, restfa1_in13_s, restfa2_in12_s, restfa2_in13_s;
  wire restfa1_in12_c, restfa1_in13_c, restfa2_in12_c, restfa2_in13_c;
  
  wire restfa1_in14_int0, restfa2_in14_int0, restfa3_in14_int0;
  wire restfa1_in14_int1, restfa2_in14_int1, restfa3_in14_int1;
  wire restfa1_in14_int2, restfa2_in14_int2, restfa3_in14_int2;
  wire restfa1_in14_s, restfa2_in14_s, restfa3_in14_s;
  wire restfa1_in14_c, restfa2_in14_c, restfa3_in14_c;

  assign n73 = ~pi06 & ~pi07;
  assign n74 = ~pi08 & n73;
  assign po00 = ~pi09 & n74;
  assign n76 = ~pi11 & ~pi12;
  assign po01 = ~pi10 | n76;
  assign n78 = pi09 & pi32;
  assign n79 = pi08 & pi31;
  assign n80 = pi06 & pi29;
  assign n81 = pi07 & pi30;
  assign n82 = ~n80 & ~n81;
  assign n83 = ~n79 & n82;
  assign n84 = ~n78 & n83;
  assign n85 = pi13 & pi36;
  assign n86 = pi12 & pi35;
  assign n87 = pi10 & pi33;
  assign n88 = pi11 & pi34;
  assign n89 = ~n87 & ~n88;
  assign n90 = ~n86 & n89;
  assign n91 = ~n85 & n90;
  assign n92 = n84 & n91;
  assign n93 = pi00 & pi01;
  assign n94 = pi02 & n93;
  assign n95 = pi00 & ~pi01;
  assign n96 = pi02 & n95;
  assign n97 = ~n94 & ~n96;
  assign n98 = ~n92 & n97;
  assign n99 = ~pi07 & ~pi08;
  assign n100 = pi06 & ~n99;
  assign n101 = n94 & n100;
  assign n102 = ~pi34 & ~pi35;
  assign n103 = pi33 & ~n102;
  assign n104 = n96 & n103;
  assign n105 = ~n101 & ~n104;
  assign po02 = ~n98 & n105;
  assign n107 = ~pi35 & pi36;
  assign n108 = pi35 & ~pi36;
  assign n109 = ~n107 & ~n108;
  assign n110 = ~pi33 & pi34;
  assign n111 = pi33 & ~pi34;
  assign n112 = ~n110 & ~n111;
  assign n113 = ~n109 & n112;
  assign n114 = n109 & ~n112;
  assign n115 = ~n113 & ~n114;
  assign n116 = ~pi31 & pi32;
  assign n117 = pi31 & ~pi32;
  assign n118 = ~n116 & ~n117;
  assign n119 = ~pi29 & pi30;
  assign n120 = pi29 & ~pi30;
  assign n121 = ~n119 & ~n120;
  assign n122 = ~n118 & n121;
  assign n123 = n118 & ~n121;
  assign n124 = ~n122 & ~n123;
  assign n125 = ~n115 & n124;
  assign n126 = n115 & ~n124;
  assign po03 = ~n125 & ~n126;
  assign n128 = pi12 & ~pi13;
  assign n129 = ~pi12 & pi13;
  assign n130 = ~n128 & ~n129;
  assign n131 = ~pi10 & ~pi11;
  assign n132 = pi10 & pi11;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~n130 & ~n133;
  assign n135 = n130 & n133;
  assign n136 = ~n134 & ~n135;
  assign n137 = pi06 & pi07;
  assign n138 = ~n73 & ~n137;
  assign n139 = pi08 & pi09;
  assign n140 = ~pi08 & ~pi09;
  assign n141 = ~n139 & ~n140;
  assign n142 = n138 & n141;
  assign n143 = ~n138 & ~n141;
  assign n144 = ~n142 & ~n143;
  assign n145 = ~n136 & n144;
  assign n146 = n136 & ~n144;
  assign po04 = n145 | n146;
  assign n148 = pi01 & pi02;
  assign n149 = ~pi00 & n148;
  assign n150 = pi03 & n96;
  assign n151 = ~n93 & ~n150;
  assign n152 = ~n149 & n151;
  assign n153 = ~pi00 & pi03;
  assign n154 = pi13 & ~n153;
  assign n155 = n152 & n154;
  assign n156 = ~pi02 & pi03;
  assign n157 = ~pi02 & ~n156;
  assign n158 = pi11 & n157;
  assign n159 = pi02 & pi13;
  assign n160 = pi38 & n156;
  assign n161 = ~n159 & ~n160;
  assign n162 = ~n158 & n161;
  assign n163 = ~n151 & ~n162;
  assign n164 = ~pi13 & n149;
  assign n165 = ~n163 & ~n164;
  assign n166 = ~n155 & n165;
  assign n167 = pi03 & pi04;
  assign n168 = n93 & ~n167;
  assign n169 = ~pi03 & ~pi48;
  assign n170 = ~pi03 & ~n169;
  assign n171 = pi35 & n170;
  assign n172 = pi03 & pi40;
  assign n173 = pi34 & n169;
  assign n174 = ~n172 & ~n173;
  assign n175 = ~n171 & n174;
  assign n176 = n168 & ~n175;
  assign n177 = pi37 & ~n168;
  assign n178 = ~pi00 & pi05;
  assign n179 = ~pi04 & n178;
  assign n180 = n177 & n179;
  assign n181 = pi36 & ~n168;
  assign n182 = ~n179 & n181;
  assign n183 = ~n180 & ~n182;
  assign n184 = ~n176 & n183;
  assign n185 = pi23 & n184;
  assign n186 = pi22 & ~n184;
  assign n187 = ~n185 & ~n186;
  assign n188 = ~n166 & ~n187;
  assign n189 = ~pi24 & n184;
  assign n190 = ~pi25 & ~n184;
  assign n191 = ~n189 & ~n190;
  assign n192 = n166 & ~n191;
  assign n193 = ~n188 & ~n192;
  assign n194 = pi12 & ~n153;
  assign n195 = n152 & n194;
  assign n196 = pi10 & n157;
  assign n197 = pi02 & ~pi12;
  assign n198 = pi13 & n156;
  assign n199 = ~n197 & ~n198;
  assign n200 = ~n196 & n199;
  assign n201 = ~n151 & ~n200;
  assign n202 = ~pi12 & n149;
  assign n203 = ~n201 & ~n202;
  assign n204 = ~n195 & n203;
  assign n205 = pi34 & n170;
  assign n206 = pi03 & pi39;
  assign n207 = pi33 & n169;
  assign n208 = ~n206 & ~n207;
  assign n209 = ~n205 & n208;
  assign n210 = n168 & ~n209;
  assign n211 = pi35 & ~n168;
  assign n212 = ~n179 & n211;
  assign n213 = ~n180 & ~n212;
  assign n214 = ~n210 & n213;
  assign n215 = pi23 & n214;
  assign n216 = pi22 & ~n214;
  assign n217 = ~n215 & ~n216;
  assign n218 = ~n204 & ~n217;
  assign n219 = ~pi24 & n214;
  assign n220 = ~pi25 & ~n214;
  assign n221 = ~n219 & ~n220;
  assign n222 = n204 & ~n221;
  assign n223 = ~n218 & ~n222;
  assign n224 = pi10 & ~n153;
  assign n225 = n152 & n224;
  assign n226 = pi08 & n157;
  assign n227 = ~pi12 & n131;
  assign n228 = pi02 & ~n227;
  assign n229 = pi11 & n156;
  assign n230 = ~n228 & ~n229;
  assign n231 = ~n226 & n230;
  assign n232 = ~n151 & ~n231;
  assign n233 = ~pi10 & n149;
  assign n234 = ~n232 & ~n233;
  assign n235 = ~n225 & n234;
  assign n236 = pi32 & n170;
  assign n237 = pi03 & pi13;
  assign n238 = pi31 & n169;
  assign n239 = ~n237 & ~n238;
  assign n240 = ~n236 & n239;
  assign n241 = n168 & ~n240;
  assign n242 = pi33 & ~n168;
  assign n243 = ~n178 & n242;
  assign n244 = n177 & n178;
  assign n245 = ~n243 & ~n244;
  assign n246 = ~n241 & n245;
  assign n247 = pi23 & n246;
  assign n248 = pi22 & ~n246;
  assign n249 = ~n247 & ~n248;
  assign n250 = ~n235 & ~n249;
  assign n251 = ~pi24 & n246;
  assign n252 = ~pi25 & ~n246;
  assign n253 = ~n251 & ~n252;
  assign n254 = n235 & ~n253;
  assign n255 = ~n250 & ~n254;
  assign n256 = pi11 & ~n153;
  assign n257 = n152 & n256;
  assign n258 = pi09 & n157;
  assign n259 = pi11 & pi12;
  assign n260 = ~n76 & ~n259;
  assign n261 = pi02 & ~n260;
  assign n262 = pi12 & n156;
  assign n263 = ~n261 & ~n262;
  assign n264 = ~n258 & n263;
  assign n265 = ~n151 & ~n264;
  assign n266 = ~pi11 & n149;
  assign n267 = ~n265 & ~n266;
  assign n268 = ~n257 & n267;
  assign n269 = pi33 & n170;
  assign n270 = pi03 & pi38;
  assign n271 = pi32 & n169;
  assign n272 = ~n270 & ~n271;
  assign n273 = ~n269 & n272;
  assign n274 = n168 & ~n273;
  assign n275 = pi34 & ~n168;
  assign n276 = ~n179 & n275;
  assign n277 = ~n180 & ~n276;
  assign n278 = ~n274 & n277;
  assign n279 = pi23 & n278;
  assign n280 = pi22 & ~n278;
  assign n281 = ~n279 & ~n280;
  assign n282 = ~n268 & ~n281;
  assign n283 = ~pi24 & n278;
  assign n284 = ~pi25 & ~n278;
  assign n285 = ~n283 & ~n284;
  assign n286 = n268 & ~n285;
  assign n287 = ~n282 & ~n286;
  assign n288 = n255 & n287;
  assign n289 = n223 & n288;
  assign n290 = n193 & n289;
  assign n291 = ~pi00 & pi02;
  assign n292 = pi09 & ~n291;
  assign n293 = n152 & n292;
  assign n294 = pi07 & n157;
  assign n295 = pi02 & pi09;
  assign n296 = pi10 & n156;
  assign n297 = ~n295 & ~n296;
  assign n298 = ~n294 & n297;
  assign n299 = ~n151 & ~n298;
  assign n300 = ~pi09 & n149;
  assign n301 = ~n299 & ~n300;
  assign n302 = ~n293 & n301;
  assign n303 = pi31 & n170;
  assign n304 = pi03 & pi12;
  assign n305 = pi30 & n169;
  assign n306 = ~n304 & ~n305;
  assign n307 = ~n303 & n306;
  assign n308 = n168 & ~n307;
  assign n309 = ~pi04 & ~pi05;
  assign n310 = ~pi00 & ~n309;
  assign n311 = n177 & n310;
  assign n312 = pi32 & ~n168;
  assign n313 = ~n310 & n312;
  assign n314 = ~n311 & ~n313;
  assign n315 = ~n308 & n314;
  assign n316 = pi23 & n315;
  assign n317 = pi22 & ~n315;
  assign n318 = ~n316 & ~n317;
  assign n319 = ~n302 & ~n318;
  assign n320 = ~pi24 & n315;
  assign n321 = ~pi25 & ~n315;
  assign n322 = ~n320 & ~n321;
  assign n323 = n302 & ~n322;
  assign n324 = ~n319 & ~n323;
  assign n325 = pi08 & ~n291;
  assign n326 = n152 & n325;
  assign n327 = pi06 & n157;
  assign n328 = pi02 & ~pi08;
  assign n329 = pi09 & n156;
  assign n330 = ~n328 & ~n329;
  assign n331 = ~n327 & n330;
  assign n332 = ~n151 & ~n331;
  assign n333 = ~pi08 & n149;
  assign n334 = ~n332 & ~n333;
  assign n335 = ~n326 & n334;
  assign n336 = pi30 & n170;
  assign n337 = pi03 & pi11;
  assign n338 = pi29 & n169;
  assign n339 = ~n337 & ~n338;
  assign n340 = ~n336 & n339;
  assign n341 = n168 & ~n340;
  assign n342 = pi31 & ~n168;
  assign n343 = ~n310 & n342;
  assign n344 = ~n311 & ~n343;
  assign n345 = ~n341 & n344;
  assign n346 = pi23 & n345;
  assign n347 = pi22 & ~n345;
  assign n348 = ~n346 & ~n347;
  assign n349 = ~n335 & ~n348;
  assign n350 = ~pi24 & n345;
  assign n351 = ~pi25 & ~n345;
  assign n352 = ~n350 & ~n351;
  assign n353 = n335 & ~n352;
  assign n354 = ~n349 & ~n353;
  assign n355 = pi06 & ~n291;
  assign n356 = n152 & n355;
  assign n357 = pi20 & n157;
  assign n358 = pi02 & ~n74;
  assign n359 = pi07 & n156;
  assign n360 = ~n358 & ~n359;
  assign n361 = ~n357 & n360;
  assign n362 = ~n151 & ~n361;
  assign n363 = ~pi06 & n149;
  assign n364 = ~n362 & ~n363;
  assign n365 = ~n356 & n364;
  assign n366 = pi28 & n170;
  assign n367 = pi03 & pi09;
  assign n368 = pi27 & n169;
  assign n369 = ~n367 & ~n368;
  assign n370 = ~n366 & n369;
  assign n371 = n168 & ~n370;
  assign n372 = pi29 & ~n168;
  assign n373 = ~n310 & n372;
  assign n374 = ~n311 & ~n373;
  assign n375 = ~n371 & n374;
  assign n376 = pi23 & n375;
  assign n377 = pi22 & ~n375;
  assign n378 = ~n376 & ~n377;
  assign n379 = ~n365 & ~n378;
  assign n380 = ~pi24 & n375;
  assign n381 = ~pi25 & ~n375;
  assign n382 = ~n380 & ~n381;
  assign n383 = n365 & ~n382;
  assign n384 = ~n379 & ~n383;
  assign n385 = pi07 & ~n291;
  assign n386 = n152 & n385;
  assign n387 = pi21 & n157;
  assign n388 = pi07 & pi08;
  assign n389 = ~n99 & ~n388;
  assign n390 = pi02 & ~n389;
  assign n391 = pi08 & n156;
  assign n392 = ~n390 & ~n391;
  assign n393 = ~n387 & n392;
  assign n394 = ~n151 & ~n393;
  assign n395 = ~pi07 & n149;
  assign n396 = ~n394 & ~n395;
  assign n397 = ~n386 & n396;
  assign n398 = pi29 & n170;
  assign n399 = pi03 & pi10;
  assign n400 = pi28 & n169;
  assign n401 = ~n399 & ~n400;
  assign n402 = ~n398 & n401;
  assign n403 = n168 & ~n402;
  assign n404 = pi30 & ~n168;
  assign n405 = ~n310 & n404;
  assign n406 = ~n311 & ~n405;
  assign n407 = ~n403 & n406;
  assign n408 = pi23 & n407;
  assign n409 = pi22 & ~n407;
  assign n410 = ~n408 & ~n409;
  assign n411 = ~n397 & ~n410;
  assign n412 = ~pi24 & n407;
  assign n413 = ~pi25 & ~n407;
  assign n414 = ~n412 & ~n413;
  assign n415 = n397 & ~n414;
  assign n416 = ~n411 & ~n415;
  assign n417 = n384 & n416;
  assign n418 = n354 & n417;
  assign n419 = n324 & n418;
  assign po05 = n290 & n419;
  assign n421 = ~n188 & ~n218;
  assign n422 = ~n222 & ~n421;
  assign n423 = ~n282 & ~n422;
  assign n424 = ~n286 & ~n423;
  assign n425 = ~n250 & ~n424;
  assign n426 = ~n254 & ~n425;
  assign n427 = n419 & n426;
  assign n428 = ~n319 & ~n349;
  assign n429 = ~n353 & ~n428;
  assign n430 = ~n411 & ~n429;
  assign n431 = ~n415 & ~n430;
  assign n432 = ~n379 & ~n431;
  assign n433 = ~n383 & ~n432;
  assign po06 = n427 | n433;
  assign n435 = ~pi00 & pi01;
  assign n436 = ~pi02 & n435;
  assign n437 = pi26 & n436;
  assign n438 = pi47 & n437;
  assign n439 = n218 & ~n438;
  assign n440 = ~n204 & n438;
  assign n441 = ~n223 & n440;
  assign n442 = n223 & ~n440;
  assign n443 = ~n441 & ~n442;
  assign n444 = n188 & ~n438;
  assign n445 = ~n443 & n444;
  assign n446 = ~n439 & ~n445;
  assign n447 = ~n166 & n438;
  assign n448 = ~n193 & n447;
  assign n449 = n193 & ~n447;
  assign n450 = ~n448 & ~n449;
  assign n451 = ~n443 & ~n450;
  assign n452 = pi46 & n451;
  assign po07 = ~n446 | n452;
  assign n454 = ~pi13 & n227;
  assign n455 = ~pi04 & n96;
  assign n456 = pi00 & ~n455;
  assign n457 = n454 & n456;
  assign n458 = n100 & n455;
  assign n459 = n426 & ~n438;
  assign n460 = ~n246 & ~n278;
  assign n461 = ~n214 & n460;
  assign n462 = ~n184 & n461;
  assign n463 = ~pi23 & n462;
  assign n464 = n246 & n278;
  assign n465 = n214 & n464;
  assign n466 = n185 & n465;
  assign n467 = ~n463 & ~n466;
  assign n468 = n438 & ~n467;
  assign n469 = n290 & ~n438;
  assign n470 = ~n468 & ~n469;
  assign n471 = pi46 & ~n470;
  assign n472 = ~n459 & ~n471;
  assign n473 = ~pi00 & ~n472;
  assign n474 = ~n458 & ~n473;
  assign po08 = n457 | ~n474;
  assign n476 = ~pi13 & ~n96;
  assign n477 = pi05 & ~n144;
  assign n478 = ~pi05 & n100;
  assign n479 = ~n477 & ~n478;
  assign n480 = n150 & n479;
  assign n481 = ~pi03 & n96;
  assign n482 = po01 & n481;
  assign n483 = ~n480 & ~n482;
  assign n484 = ~n476 & n483;
  assign n485 = pi02 & ~pi22;
  assign n486 = n93 & ~n485;
  assign n487 = ~pi01 & ~pi02;
  assign n488 = ~pi03 & n487;
  assign n489 = ~n486 & ~n488;
  assign n490 = ~n484 & n489;
  assign n491 = pi02 & ~pi24;
  assign n492 = pi02 & pi23;
  assign n493 = pi25 & n492;
  assign n494 = ~n491 & n493;
  assign n495 = pi06 & n494;
  assign n496 = ~pi25 & n492;
  assign n497 = ~n491 & n496;
  assign n498 = pi07 & n497;
  assign n499 = n491 & n493;
  assign n500 = pi08 & n499;
  assign n501 = n491 & n496;
  assign n502 = pi09 & n501;
  assign n503 = pi02 & pi25;
  assign n504 = ~n492 & n503;
  assign n505 = ~n491 & n504;
  assign n506 = pi10 & n505;
  assign n507 = ~n492 & ~n503;
  assign n508 = ~n491 & n507;
  assign n509 = pi11 & n508;
  assign n510 = n491 & n507;
  assign n511 = pi21 & n510;
  assign n512 = n491 & n504;
  assign n513 = pi12 & n512;
  assign n514 = ~n511 & ~n513;
  assign n515 = ~n509 & n514;
  assign n516 = ~n506 & n515;
  assign n517 = ~n502 & n516;
  assign n518 = ~n500 & n517;
  assign n519 = ~n498 & n518;
  assign n520 = ~n495 & n519;
  assign n521 = ~pi03 & n520;
  assign n522 = pi44 & n494;
  assign n523 = pi43 & n497;
  assign n524 = pi42 & n499;
  assign n525 = pi41 & n501;
  assign n526 = pi40 & n505;
  assign n527 = pi39 & n508;
  assign n528 = pi45 & n510;
  assign n529 = pi38 & n512;
  assign n530 = ~n528 & ~n529;
  assign n531 = ~n527 & n530;
  assign n532 = ~n526 & n531;
  assign n533 = ~n525 & n532;
  assign n534 = ~n524 & n533;
  assign n535 = ~n523 & n534;
  assign n536 = ~n522 & n535;
  assign n537 = pi03 & n536;
  assign n538 = ~n521 & ~n537;
  assign n539 = n486 & ~n538;
  assign n540 = n450 & n488;
  assign n541 = ~n539 & ~n540;
  assign n542 = ~n490 & n541;
  assign n543 = pi01 & ~pi02;
  assign n544 = pi05 & n543;
  assign n545 = pi00 & ~n544;
  assign n546 = ~n455 & n545;
  assign n547 = n542 & n546;
  assign n548 = pi46 & ~n450;
  assign n549 = ~pi46 & n450;
  assign n550 = ~n546 & ~n549;
  assign n551 = ~n548 & n550;
  assign po09 = n547 | n551;
  assign n553 = ~pi01 & ~pi03;
  assign n554 = ~n486 & ~n553;
  assign n555 = ~pi09 & n554;
  assign n556 = pi18 & n494;
  assign n557 = pi19 & n497;
  assign n558 = pi20 & n499;
  assign n559 = pi21 & n501;
  assign n560 = pi06 & n505;
  assign n561 = pi07 & n508;
  assign n562 = pi17 & n510;
  assign n563 = pi08 & n512;
  assign n564 = ~n562 & ~n563;
  assign n565 = ~n561 & n564;
  assign n566 = ~n560 & n565;
  assign n567 = ~n559 & n566;
  assign n568 = ~n558 & n567;
  assign n569 = ~n557 & n568;
  assign n570 = ~n556 & n569;
  assign n571 = ~pi03 & n570;
  assign n572 = pi40 & n494;
  assign n573 = pi39 & n497;
  assign n574 = pi38 & n499;
  assign n575 = pi13 & n501;
  assign n576 = pi12 & n505;
  assign n577 = pi41 & n510;
  assign n578 = pi10 & n512;
  assign n579 = ~n577 & ~n578;
  assign n580 = ~n509 & n579;
  assign n581 = ~n576 & n580;
  assign n582 = ~n575 & n581;
  assign n583 = ~n574 & n582;
  assign n584 = ~n573 & n583;
  assign n585 = ~n572 & n584;
  assign n586 = pi03 & n585;
  assign n587 = ~n571 & ~n586;
  assign n588 = n486 & ~n587;
  assign n589 = ~n302 & n438;
  assign n590 = ~n324 & n589;
  assign n591 = n324 & ~n589;
  assign n592 = ~n590 & ~n591;
  assign n593 = n553 & n592;
  assign n594 = ~n588 & ~n593;
  assign n595 = ~n555 & n594;
  assign n596 = n546 & n595;
  assign n597 = n459 & ~n592;
  assign n598 = ~n459 & n592;
  assign n599 = ~n597 & ~n598;
  assign n600 = n471 & ~n599;
  assign n601 = ~n471 & n599;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~n545 & ~n602;
  assign n604 = n455 & ~n602;
  assign n605 = ~n603 & ~n604;
  assign po10 = n596 | ~n605;
  assign n607 = n419 & ~n470;
  assign n608 = ~n397 & n437;
  assign n609 = ~n416 & n608;
  assign n610 = n416 & ~n608;
  assign n611 = ~n609 & ~n610;
  assign n612 = ~n470 & ~n611;
  assign n613 = ~n335 & n438;
  assign n614 = ~n354 & n613;
  assign n615 = n354 & ~n613;
  assign n616 = ~n614 & ~n615;
  assign n617 = ~n592 & ~n616;
  assign n618 = n612 & n617;
  assign n619 = ~n607 & n618;
  assign n620 = n607 & ~n618;
  assign n621 = ~n619 & ~n620;
  assign n622 = pi46 & ~n621;
  assign n623 = n419 & n459;
  assign n624 = ~n433 & ~n623;
  assign n625 = ~n611 & ~n616;
  assign n626 = n319 & ~n438;
  assign n627 = n625 & n626;
  assign n628 = n411 & ~n437;
  assign n629 = n349 & ~n438;
  assign n630 = ~n611 & n629;
  assign n631 = ~n628 & ~n630;
  assign n632 = ~n627 & n631;
  assign n633 = n597 & n625;
  assign n634 = n632 & ~n633;
  assign n635 = ~n624 & n634;
  assign n636 = n624 & ~n634;
  assign n637 = ~n635 & ~n636;
  assign n638 = n622 & n637;
  assign n639 = ~n622 & ~n637;
  assign n640 = ~n638 & ~n639;
  assign n641 = ~n94 & ~n95;
  assign n642 = ~n640 & n641;
  assign n643 = pi09 & n389;
  assign n644 = pi06 & n643;
  assign n645 = ~pi06 & pi08;
  assign n646 = ~n644 & ~n645;
  assign n647 = n95 & ~n646;
  assign n648 = pi13 & n260;
  assign n649 = n94 & n648;
  assign n650 = ~n647 & ~n649;
  assign po11_prelocked = n642 | ~n650;
  assign n652 = n115 & n150;
  assign n653 = pi10 & ~n96;
  assign n654 = ~n652 & ~n653;
  assign n655 = n489 & n654;
  assign n656 = pi19 & n494;
  assign n657 = pi20 & n497;
  assign n658 = pi21 & n499;
  assign n659 = pi06 & n501;
  assign n660 = pi07 & n505;
  assign n661 = pi08 & n508;
  assign n662 = pi18 & n510;
  assign n663 = pi09 & n512;
  assign n664 = ~n662 & ~n663;
  assign n665 = ~n661 & n664;
  assign n666 = ~n660 & n665;
  assign n667 = ~n659 & n666;
  assign n668 = ~n658 & n667;
  assign n669 = ~n657 & n668;
  assign n670 = ~n656 & n669;
  assign n671 = ~pi03 & n670;
  assign n672 = pi41 & n494;
  assign n673 = pi40 & n497;
  assign n674 = pi39 & n499;
  assign n675 = pi38 & n501;
  assign n676 = pi13 & n505;
  assign n677 = pi12 & n508;
  assign n678 = pi42 & n510;
  assign n679 = pi11 & n512;
  assign n680 = ~n678 & ~n679;
  assign n681 = ~n677 & n680;
  assign n682 = ~n676 & n681;
  assign n683 = ~n675 & n682;
  assign n684 = ~n674 & n683;
  assign n685 = ~n673 & n684;
  assign n686 = ~n672 & n685;
  assign n687 = pi03 & n686;
  assign n688 = ~n671 & ~n687;
  assign n689 = n486 & ~n688;
  assign n690 = ~n235 & n438;
  assign n691 = ~n255 & n690;
  assign n692 = n255 & ~n690;
  assign n693 = ~n691 & ~n692;
  assign n694 = n488 & n693;
  assign n695 = ~n689 & ~n694;
  assign n696 = ~n655 & n695;
  assign n697 = n546 & n696;
  assign n698 = ~n268 & n438;
  assign n699 = ~n287 & n698;
  assign n700 = n287 & ~n698;
  assign n701 = ~n699 & ~n700;
  assign n702 = n451 & ~n701;
  assign n703 = pi46 & n702;
  assign n704 = n188 & ~n443;
  assign n705 = ~n218 & ~n704;
  assign n706 = ~n701 & ~n705;
  assign n707 = ~n282 & ~n706;
  assign n708 = ~n438 & ~n707;
  assign n709 = ~n693 & ~n708;
  assign n710 = n693 & n708;
  assign n711 = ~n709 & ~n710;
  assign n712 = n703 & n711;
  assign n713 = ~n703 & ~n711;
  assign n714 = ~n712 & ~n713;
  assign n715 = ~n545 & ~n714;
  assign n716 = n443 & ~n444;
  assign n717 = ~n445 & ~n716;
  assign n718 = n548 & ~n717;
  assign n719 = ~n548 & n717;
  assign n720 = ~n718 & ~n719;
  assign n721 = n446 & ~n701;
  assign n722 = ~n446 & n701;
  assign n723 = ~n721 & ~n722;
  assign n724 = n452 & n723;
  assign n725 = ~n452 & ~n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = ~n720 & ~n726;
  assign n728 = n472 & ~n727;
  assign n729 = ~n714 & ~n728;
  assign n730 = n455 & n729;
  assign n731 = ~n715 & ~n730;
  assign po12_prelocked = n697 | ~n731;
  assign n733 = ~pi12 & ~n96;
  assign n734 = pi05 & n124;
  assign n735 = ~n139 & n454;
  assign n736 = ~pi06 & n735;
  assign n737 = pi07 & n736;
  assign n738 = ~pi05 & n737;
  assign n739 = ~n734 & ~n738;
  assign n740 = n150 & n739;
  assign n741 = ~n454 & n481;
  assign n742 = ~n740 & ~n741;
  assign n743 = ~n733 & n742;
  assign n744 = n489 & ~n743;
  assign n745 = pi21 & n494;
  assign n746 = pi06 & n497;
  assign n747 = pi07 & n499;
  assign n748 = pi08 & n501;
  assign n749 = pi09 & n505;
  assign n750 = pi10 & n508;
  assign n751 = pi20 & n510;
  assign n752 = ~n679 & ~n751;
  assign n753 = ~n750 & n752;
  assign n754 = ~n749 & n753;
  assign n755 = ~n748 & n754;
  assign n756 = ~n747 & n755;
  assign n757 = ~n746 & n756;
  assign n758 = ~n745 & n757;
  assign n759 = ~pi03 & n758;
  assign n760 = pi43 & n494;
  assign n761 = pi42 & n497;
  assign n762 = pi41 & n499;
  assign n763 = pi40 & n501;
  assign n764 = pi39 & n505;
  assign n765 = pi38 & n508;
  assign n766 = pi44 & n510;
  assign n767 = pi13 & n512;
  assign n768 = ~n766 & ~n767;
  assign n769 = ~n765 & n768;
  assign n770 = ~n764 & n769;
  assign n771 = ~n763 & n770;
  assign n772 = ~n762 & n771;
  assign n773 = ~n761 & n772;
  assign n774 = ~n760 & n773;
  assign n775 = pi03 & n774;
  assign n776 = ~n759 & ~n775;
  assign n777 = n486 & ~n776;
  assign n778 = n443 & n488;
  assign n779 = ~n777 & ~n778;
  assign n780 = ~n744 & n779;
  assign n781 = n546 & n780;
  assign n782 = ~n545 & ~n720;
  assign n783 = n472 & ~n720;
  assign n784 = ~n472 & n720;
  assign n785 = ~n783 & ~n784;
  assign n786 = n455 & n785;
  assign n787 = ~n782 & ~n786;
  assign po13_prelocked = n781 | ~n787;
  assign n789 = n136 & n150;
  assign n790 = pi11 & ~n96;
  assign n791 = ~n789 & ~n790;
  assign n792 = n489 & n791;
  assign n793 = pi20 & n494;
  assign n794 = pi21 & n497;
  assign n795 = pi06 & n499;
  assign n796 = pi07 & n501;
  assign n797 = pi08 & n505;
  assign n798 = pi09 & n508;
  assign n799 = pi19 & n510;
  assign n800 = ~n578 & ~n799;
  assign n801 = ~n798 & n800;
  assign n802 = ~n797 & n801;
  assign n803 = ~n796 & n802;
  assign n804 = ~n795 & n803;
  assign n805 = ~n794 & n804;
  assign n806 = ~n793 & n805;
  assign n807 = ~pi03 & n806;
  assign n808 = pi42 & n494;
  assign n809 = pi41 & n497;
  assign n810 = pi40 & n499;
  assign n811 = pi39 & n501;
  assign n812 = pi38 & n505;
  assign n813 = pi13 & n508;
  assign n814 = pi43 & n510;
  assign n815 = ~n513 & ~n814;
  assign n816 = ~n813 & n815;
  assign n817 = ~n812 & n816;
  assign n818 = ~n811 & n817;
  assign n819 = ~n810 & n818;
  assign n820 = ~n809 & n819;
  assign n821 = ~n808 & n820;
  assign n822 = pi03 & n821;
  assign n823 = ~n807 & ~n822;
  assign n824 = n486 & ~n823;
  assign n825 = n488 & n701;
  assign n826 = ~n824 & ~n825;
  assign n827 = ~n792 & n826;
  assign n828 = n546 & n827;
  assign n829 = ~n545 & ~n726;
  assign n830 = n726 & n783;
  assign n831 = ~n726 & ~n783;
  assign n832 = ~n830 & ~n831;
  assign n833 = n455 & ~n832;
  assign n834 = ~n829 & ~n833;
  assign po14_prelocked = n828 | ~n834;
  assign n836 = ~pi07 & n554;
  assign n837 = pi16 & n494;
  assign n838 = pi17 & n497;
  assign n839 = pi18 & n499;
  assign n840 = pi19 & n501;
  assign n841 = pi20 & n505;
  assign n842 = pi21 & n508;
  assign n843 = pi15 & n510;
  assign n844 = pi06 & n512;
  assign n845 = ~n843 & ~n844;
  assign n846 = ~n842 & n845;
  assign n847 = ~n841 & n846;
  assign n848 = ~n840 & n847;
  assign n849 = ~n839 & n848;
  assign n850 = ~n838 & n849;
  assign n851 = ~n837 & n850;
  assign n852 = ~pi03 & n851;
  assign n853 = pi38 & n494;
  assign n854 = pi13 & n497;
  assign n855 = pi12 & n499;
  assign n856 = pi11 & n501;
  assign n857 = pi39 & n510;
  assign n858 = ~n563 & ~n857;
  assign n859 = ~n798 & n858;
  assign n860 = ~n506 & n859;
  assign n861 = ~n856 & n860;
  assign n862 = ~n855 & n861;
  assign n863 = ~n854 & n862;
  assign n864 = ~n853 & n863;
  assign n865 = pi03 & n864;
  assign n866 = ~n852 & ~n865;
  assign n867 = n486 & ~n866;
  assign n868 = n553 & n611;
  assign n869 = ~n867 & ~n868;
  assign n870 = ~n836 & n869;
  assign n871 = n546 & n870;
  assign n872 = ~n470 & ~n592;
  assign n873 = ~n616 & n872;
  assign n874 = pi46 & n873;
  assign n875 = n459 & n617;
  assign n876 = ~n616 & n626;
  assign n877 = ~n629 & ~n876;
  assign n878 = ~n875 & n877;
  assign n879 = ~n611 & n878;
  assign n880 = n611 & ~n878;
  assign n881 = ~n879 & ~n880;
  assign n882 = n874 & n881;
  assign n883 = ~n874 & ~n881;
  assign n884 = ~n882 & ~n883;
  assign n885 = ~n545 & ~n884;
  assign n886 = pi46 & n872;
  assign n887 = ~n597 & ~n626;
  assign n888 = ~n616 & n887;
  assign n889 = n616 & ~n887;
  assign n890 = ~n888 & ~n889;
  assign n891 = n886 & n890;
  assign n892 = ~n886 & ~n890;
  assign n893 = ~n891 & ~n892;
  assign n894 = pi46 & n607;
  assign n895 = n624 & ~n894;
  assign n896 = ~n893 & n895;
  assign n897 = n884 & n896;
  assign n898 = ~n884 & ~n896;
  assign n899 = ~n897 & ~n898;
  assign n900 = n455 & ~n899;
  assign n901 = ~n885 & ~n900;
  assign po15_prelocked = n871 | ~n901;
  assign n903 = ~pi06 & n554;
  assign n904 = pi04 & ~pi06;
  assign n905 = ~pi03 & ~pi04;
  assign n906 = pi15 & n494;
  assign n907 = pi16 & n497;
  assign n908 = pi17 & n499;
  assign n909 = pi18 & n501;
  assign n910 = pi19 & n505;
  assign n911 = pi20 & n508;
  assign n912 = pi14 & n510;
  assign n913 = pi21 & n512;
  assign n914 = ~n912 & ~n913;
  assign n915 = ~n911 & n914;
  assign n916 = ~n910 & n915;
  assign n917 = ~n909 & n916;
  assign n918 = ~n908 & n917;
  assign n919 = ~n907 & n918;
  assign n920 = ~n906 & n919;
  assign n921 = n905 & n920;
  assign n922 = pi03 & ~pi04;
  assign n923 = pi13 & n494;
  assign n924 = pi12 & n497;
  assign n925 = pi11 & n499;
  assign n926 = pi10 & n501;
  assign n927 = pi38 & n510;
  assign n928 = pi07 & n512;
  assign n929 = ~n927 & ~n928;
  assign n930 = ~n661 & n929;
  assign n931 = ~n749 & n930;
  assign n932 = ~n926 & n931;
  assign n933 = ~n925 & n932;
  assign n934 = ~n924 & n933;
  assign n935 = ~n923 & n934;
  assign n936 = n922 & n935;
  assign n937 = ~n921 & ~n936;
  assign n938 = ~n904 & n937;
  assign n939 = n486 & ~n938;
  assign n940 = ~n365 & n437;
  assign n941 = ~n384 & n940;
  assign n942 = n384 & ~n940;
  assign n943 = ~n941 & ~n942;
  assign n944 = n553 & n943;
  assign n945 = ~n939 & ~n944;
  assign n946 = ~n903 & n945;
  assign n947 = n546 & n946;
  assign n948 = pi46 & n618;
  assign n949 = n634 & ~n943;
  assign n950 = ~n634 & n943;
  assign n951 = ~n949 & ~n950;
  assign n952 = n948 & n951;
  assign n953 = ~n948 & ~n951;
  assign n954 = ~n952 & ~n953;
  assign n955 = ~n545 & ~n954;
  assign n956 = ~n884 & ~n893;
  assign n957 = n895 & ~n956;
  assign n958 = ~n954 & ~n957;
  assign n959 = n455 & n958;
  assign n960 = ~n955 & ~n959;
  assign po16_prelocked = n947 | ~n960;
  assign n962 = ~pi08 & n554;
  assign n963 = pi17 & n494;
  assign n964 = pi18 & n497;
  assign n965 = pi19 & n499;
  assign n966 = pi20 & n501;
  assign n967 = pi21 & n505;
  assign n968 = pi06 & n508;
  assign n969 = pi16 & n510;
  assign n970 = ~n928 & ~n969;
  assign n971 = ~n968 & n970;
  assign n972 = ~n967 & n971;
  assign n973 = ~n966 & n972;
  assign n974 = ~n965 & n973;
  assign n975 = ~n964 & n974;
  assign n976 = ~n963 & n975;
  assign n977 = ~pi03 & n976;
  assign n978 = pi39 & n494;
  assign n979 = pi38 & n497;
  assign n980 = pi13 & n499;
  assign n981 = pi12 & n501;
  assign n982 = pi11 & n505;
  assign n983 = pi40 & n510;
  assign n984 = ~n663 & ~n983;
  assign n985 = ~n750 & n984;
  assign n986 = ~n982 & n985;
  assign n987 = ~n981 & n986;
  assign n988 = ~n980 & n987;
  assign n989 = ~n979 & n988;
  assign n990 = ~n978 & n989;
  assign n991 = pi03 & n990;
  assign n992 = ~n977 & ~n991;
  assign n993 = n486 & ~n992;
  assign n994 = n553 & n616;
  assign n995 = ~n993 & ~n994;
  assign n996 = ~n962 & n995;
  assign n997 = n546 & n996;
  assign n998 = ~n545 & ~n893;
  assign n999 = n893 & ~n895;
  assign n1000 = ~n896 & ~n999;
  assign n1001 = n455 & n1000;
  assign n1002 = ~n998 & ~n1001;
  assign po17_prelocked = n997 | ~n1002;
  assign n1004 = ~po09 & ~po13_prelocked;
  assign n1005 = ~po14_prelocked & n1004;
  assign n1006 = ~po12_prelocked & n1005;
  assign n1007 = ~po10 & ~po17_prelocked;
  assign n1008 = ~po15_prelocked & ~po16_prelocked;
  assign n1009 = n1007 & n1008;
  assign po18_prelocked = ~n1006 | ~n1009;
  assign n1011 = pi26 & ~pi47;
  assign n1012 = n1008 & n1011;
  assign n1013 = po18_prelocked & ~n1012;
  assign po19_prelocked = ~pi26 | ~n1013;
  assign n1015 = po12_prelocked & ~po14_prelocked;
  assign n1016 = ~po12_prelocked & po14_prelocked;
  assign n1017 = ~n1015 & ~n1016;
  assign n1018 = po09 & po13_prelocked;
  assign n1019 = ~n1004 & ~n1018;
  assign n1020 = ~n1017 & ~n1019;
  assign n1021 = n1017 & n1019;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = po10 & po17_prelocked;
  assign n1024 = ~n1007 & ~n1023;
  assign n1025 = po15_prelocked & po16_prelocked;
  assign n1026 = ~n1008 & ~n1025;
  assign n1027 = ~n1011 & n1026;
  assign n1028 = ~n1024 & n1027;
  assign n1029 = pi49 & n1011;
  assign n1030 = n1024 & ~n1027;
  assign n1031 = ~n1029 & n1030;
  assign n1032 = ~n1028 & ~n1031;
  assign n1033 = ~n1024 & n1029;
  assign n1034 = n1032 & ~n1033;
  assign n1035 = n1022 & n1034;
  assign n1036 = ~n1022 & ~n1034;
  assign po20_prelocked = n1035 | n1036;
  assign n1038 = ~n1024 & n1026;
  assign n1039 = n1024 & ~n1026;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = n1022 & ~n1040;
  assign n1042 = ~n1022 & n1040;
  assign po21_prelocked = ~n1041 & ~n1042;
  




  assign sp_in0 = n1041;
  assign sp_in1 = n115;
  assign sp_in2 = n87;
  assign sp_in3 = n642;
  assign sp_in4 = n1035;
  assign sp_in5 = n731;
  assign sp_in6 = n1004;
  assign sp_in7 = n809;
  assign sp_in8 = n781;
  assign sp_in9 = n828;
  assign sp_in10 = n901;
  assign sp_in11 = n170;
  assign sp_in12 = n960;
  assign sp_in13 = n1002;
  assign sp_in14 = n319;
  assign sp_in15 = pi26;



  assign sp_sf_in0 = sp_in0^1'b0;
  assign sp_sf_in1 = sp_in1^1'b1;
  assign sp_sf_in2 = sp_in2^1'b0;
  assign sp_sf_in3 = sp_in3^1'b0;
  assign sp_sf_in4 = sp_in4^1'b1;
  assign sp_sf_in5 = sp_in5^1'b0;
  assign sp_sf_in6 = sp_in6^1'b1;
  assign sp_sf_in7 = sp_in7^1'b0;
  assign sp_sf_in8 = sp_in8^1'b0;
  assign sp_sf_in9 = sp_in9^1'b1;
  assign sp_sf_in10 = sp_in10^1'b1;
  assign sp_sf_in11 = sp_in11^1'b1;
  assign sp_sf_in12 = sp_in12^1'b0;
  assign sp_sf_in13 = sp_in13^1'b0;
  assign sp_sf_in14 = sp_in14^1'b0;
  assign sp_sf_in15 = sp_in15^1'b1;


  assign sf_in0_s = sp_sf_in0 ^ sp_sf_in1;
  assign sf_in0_c = sp_sf_in0 & sp_sf_in1;
  assign sf_in1_s = sp_sf_in2 ^ sp_sf_in3;
  assign sf_in1_c = sp_sf_in2 & sp_sf_in3;
  assign sf_in2_s = sp_sf_in4 ^ sp_sf_in5;
  assign sf_in2_c = sp_sf_in4 & sp_sf_in5;
  assign sf_in3_s = sp_sf_in6 ^ sp_sf_in7;
  assign sf_in3_c = sp_sf_in6 & sp_sf_in7;
  assign sf_in4_s = sp_sf_in8 ^ sp_sf_in9;
  assign sf_in4_c = sp_sf_in8 & sp_sf_in9;
  assign sf_in5_s = sp_sf_in10 ^ sp_sf_in11;
  assign sf_in5_c = sp_sf_in10 & sp_sf_in11;
  assign sf_in6_s = sp_sf_in12 ^ sp_sf_in13;
  assign sf_in6_c = sp_sf_in12 & sp_sf_in13;
  assign sf_in7_s = sp_sf_in14 ^ sp_sf_in15;
  assign sf_in7_c = sp_sf_in14 & sp_sf_in15;



  assign sf_in8_s = sf_in0_s ^ sf_in1_s;
  assign sf_in8_c = sf_in0_s & sf_in1_s;
  assign fa_in8_int0 = sf_in0_c ^ sf_in1_c;
  assign fa_in8_int1 = sf_in0_c & sf_in1_c;
  assign fa_in8_int2 = sf_in8_c & fa_in8_int0;
  assign fa_in8_s = fa_in8_int0 ^ sf_in8_c;
  assign fa_in8_c = fa_in8_int1 | fa_in8_int2;

  assign sf_in9_s = sf_in2_s ^ sf_in3_s;
  assign sf_in9_c = sf_in2_s & sf_in3_s;
  assign fa_in9_int0 = sf_in2_c ^ sf_in3_c;
  assign fa_in9_int1 = sf_in2_c & sf_in3_c;
  assign fa_in9_int2 = sf_in9_c & fa_in9_int0;
  assign fa_in9_s = fa_in9_int0 ^ sf_in9_c;
  assign fa_in9_c = fa_in9_int1 | fa_in9_int2;

  assign sf_in10_s = sf_in4_s ^ sf_in5_s;
  assign sf_in10_c = sf_in4_s & sf_in5_s;
  assign fa_in10_int0 = sf_in4_c ^ sf_in5_c;
  assign fa_in10_int1 = sf_in4_c & sf_in5_c;
  assign fa_in10_int2 = sf_in10_c & fa_in10_int0;
  assign fa_in10_s = fa_in10_int0 ^ sf_in10_c;
  assign fa_in10_c = fa_in10_int1 | fa_in10_int2;

  assign sf_in11_s = sf_in6_s ^ sf_in7_s;
  assign sf_in11_c = sf_in6_s & sf_in7_s;
  assign fa_in11_int0 = sf_in6_c ^ sf_in7_c;
  assign fa_in11_int1 = sf_in6_c & sf_in7_c;
  assign fa_in11_int2 = sf_in11_c & fa_in11_int0;
  assign fa_in11_s = fa_in11_int0 ^ sf_in11_c;
  assign fa_in11_c = fa_in11_int1 | fa_in11_int2;






  assign sf_in12_s = sf_in8_s ^ sf_in9_s;
  assign sf_in12_c = sf_in8_s & sf_in9_s;
  assign fa1_in12_int0 = fa_in8_s ^ fa_in9_s;
  assign fa1_in12_int1 = fa_in8_s & fa_in9_s;
  assign fa1_in12_int2 = sf_in12_c & fa1_in12_int0;
  assign fa1_in12_s = fa1_in12_int0 ^ sf_in12_c;
  assign fa1_in12_c = fa1_in12_int1 | fa1_in12_int2;
  assign fa2_in12_int0 = fa_in8_c ^ fa_in9_c;
  assign fa2_in12_int1 = fa_in8_c & fa_in9_c;
  assign fa2_in12_int2 = fa1_in12_c & fa2_in12_int0;
  assign fa2_in12_s = fa2_in12_int0 ^ fa1_in12_c;
  assign fa2_in12_c = fa2_in12_int1 | fa2_in12_int2;
  
  assign sf_in13_s = sf_in10_s ^ sf_in11_s;
  assign sf_in13_c = sf_in10_s & sf_in11_s;
  assign fa1_in13_int0 = fa_in10_s ^ fa_in11_s;
  assign fa1_in13_int1 = fa_in10_s & fa_in11_s;
  assign fa1_in13_int2 = sf_in13_c & fa1_in13_int0;
  assign fa1_in13_s = fa1_in13_int0 ^ sf_in13_c;
  assign fa1_in13_c = fa1_in13_int1 | fa1_in13_int2;
  assign fa2_in13_int0 = fa_in10_c ^ fa_in11_c;
  assign fa2_in13_int1 = fa_in10_c & fa_in11_c;
  assign fa2_in13_int2 = fa1_in13_c & fa2_in13_int0;
  assign fa2_in13_s = fa2_in13_int0 ^ fa1_in13_c;
  assign fa2_in13_c = fa2_in13_int1 | fa2_in13_int2;
  
  



   
  
  assign sf_in14_s = sf_in12_s ^ sf_in13_s;
  assign sf_in14_c = sf_in12_s & sf_in13_s;
  assign fa1_in14_int0 = fa1_in12_s ^ fa1_in13_s;
  assign fa1_in14_int1 = fa1_in12_s & fa1_in13_s;
  assign fa1_in14_int2 = sf_in14_c & fa1_in14_int0;
  assign fa1_in14_s = fa1_in14_int0 ^ sf_in14_c;
  assign fa1_in14_c = fa1_in14_int1 | fa1_in14_int2;
  assign fa2_in14_int0 = fa2_in12_s ^ fa2_in13_s;
  assign fa2_in14_int1 = fa2_in12_s & fa2_in13_s;
  assign fa2_in14_int2 = fa1_in14_c & fa2_in14_int0;
  assign fa2_in14_s = fa2_in14_int0 ^ fa1_in14_c;
  assign fa2_in14_c = fa2_in14_int1 | fa2_in14_int2;
  assign fa3_in14_int0 = fa2_in12_c ^ fa2_in13_c;
  assign fa3_in14_int1 = fa2_in12_c & fa2_in13_c;
  assign fa3_in14_int2 = fa2_in14_c & fa3_in14_int0;
  assign fa3_in14_s = fa3_in14_int0 ^ fa2_in14_c;
  assign fa3_in14_c = fa3_in14_int1 | fa3_in14_int2;



  assign hd = (~fa3_in14_c) & (~fa3_in14_s) & (~fa2_in14_s) & (~fa1_in14_s) & sf_in14_s;
  //assign hd = (~fa3_in14_c) & (~fa3_in14_s) & (~fa2_in14_s) & (fa1_in14_s) & (~sf_in14_s);
  //assign hd = (~fa3_in14_c) & (~fa3_in14_s) & (~fa2_in14_s) & (fa1_in14_s) & sf_in14_s;


  assign rest0 = sp_in0^keyinput0;
  assign rest1 = sp_in1^keyinput1;
  assign rest2 = sp_in2^keyinput2;
  assign rest3 = sp_in3^keyinput3;
  assign rest4 = sp_in4^keyinput4;
  assign rest5 = sp_in5^keyinput5;
  assign rest6 = sp_in6^keyinput6;
  assign rest7 = sp_in7^keyinput7;
  assign rest8 = sp_in8^keyinput8;
  assign rest9 = sp_in9^keyinput9;
  assign rest10 = sp_in10^keyinput10;
  assign rest11 = sp_in11^keyinput11;
  assign rest12 = sp_in12^keyinput12;
  assign rest13 = sp_in13^keyinput13;
  assign rest14 = sp_in14^keyinput14;
  assign rest15 = sp_in15^keyinput15;

  assign rest_in0_s = rest0 ^ rest1;
  assign rest_in0_c = rest0 & rest1;
  assign rest_in1_s = rest2 ^ rest3;
  assign rest_in1_c = rest2 & rest3;
  assign rest_in2_s = rest4 ^ rest5;
  assign rest_in2_c = rest4 & rest5;
  assign rest_in3_s = rest6 ^ rest7;
  assign rest_in3_c = rest6 & rest7;
  assign rest_in4_s = rest8 ^ rest9;
  assign rest_in4_c = rest8 & rest9;
  assign rest_in5_s = rest10 ^ rest11;
  assign rest_in5_c = rest10 & rest11;
  assign rest_in6_s = rest12 ^ rest13;
  assign rest_in6_c = rest12 & rest13;
  assign rest_in7_s = rest14 ^ rest15;
  assign rest_in7_c = rest14 & rest15;

  assign rest_in8_s = rest_in0_s ^ rest_in1_s;
  assign rest_in8_c = rest_in0_s & rest_in1_s;
  assign restfa_in8_int0 = rest_in0_c ^ rest_in1_c;
  assign restfa_in8_int1 = rest_in0_c & rest_in1_c;
  assign restfa_in8_int2 = rest_in8_c & restfa_in8_int0;
  assign restfa_in8_s = restfa_in8_int0 ^ rest_in8_c;
  assign restfa_in8_c = restfa_in8_int1 | restfa_in8_int2;

  assign rest_in9_s = rest_in2_s ^ rest_in3_s;
  assign rest_in9_c = rest_in2_s & rest_in3_s;
  assign restfa_in9_int0 = rest_in2_c ^ rest_in3_c;
  assign restfa_in9_int1 = rest_in2_c & rest_in3_c;
  assign restfa_in9_int2 = rest_in9_c & restfa_in9_int0;
  assign restfa_in9_s = restfa_in9_int0 ^ rest_in9_c;
  assign restfa_in9_c = restfa_in9_int1 | restfa_in9_int2;

  assign rest_in10_s = rest_in4_s ^ rest_in5_s;
  assign rest_in10_c = rest_in4_s & rest_in5_s;
  assign restfa_in10_int0 = rest_in4_c ^ rest_in5_c;
  assign restfa_in10_int1 = rest_in4_c & rest_in5_c;
  assign restfa_in10_int2 = rest_in10_c & restfa_in10_int0;
  assign restfa_in10_s = restfa_in10_int0 ^ rest_in10_c;
  assign restfa_in10_c = restfa_in10_int1 | restfa_in10_int2;

  assign rest_in11_s = rest_in6_s ^ rest_in7_s;
  assign rest_in11_c = rest_in6_s & rest_in7_s;
  assign restfa_in11_int0 = rest_in6_c ^ rest_in7_c;
  assign restfa_in11_int1 = rest_in6_c & rest_in7_c;
  assign restfa_in11_int2 = rest_in11_c & restfa_in11_int0;
  assign restfa_in11_s = restfa_in11_int0 ^ rest_in11_c;
  assign restfa_in11_c = restfa_in11_int1 | restfa_in11_int2;







  assign rest_in12_s = rest_in8_s ^ rest_in9_s;
  assign rest_in12_c = rest_in8_s & rest_in9_s;
  assign restfa1_in12_int0 = restfa_in8_s ^ restfa_in9_s;
  assign restfa1_in12_int1 = restfa_in8_s & restfa_in9_s;
  assign restfa1_in12_int2 = rest_in12_c & restfa1_in12_int0;
  assign restfa1_in12_s = restfa1_in12_int0 ^ rest_in12_c;
  assign restfa1_in12_c = restfa1_in12_int1 | restfa1_in12_int2;
  assign restfa2_in12_int0 = restfa_in8_c ^ restfa_in9_c;
  assign restfa2_in12_int1 = restfa_in8_c & restfa_in9_c;
  assign restfa2_in12_int2 = restfa1_in12_c & restfa2_in12_int0;
  assign restfa2_in12_s = restfa2_in12_int0 ^ restfa1_in12_c;
  assign restfa2_in12_c = restfa2_in12_int1 | restfa2_in12_int2;
  
  assign rest_in13_s = rest_in10_s ^ rest_in11_s;
  assign rest_in13_c = rest_in10_s & rest_in11_s;
  assign restfa1_in13_int0 = restfa_in10_s ^ restfa_in11_s;
  assign restfa1_in13_int1 = restfa_in10_s & restfa_in11_s;
  assign restfa1_in13_int2 = rest_in13_c & restfa1_in13_int0;
  assign restfa1_in13_s = restfa1_in13_int0 ^ rest_in13_c;
  assign restfa1_in13_c = restfa1_in13_int1 | restfa1_in13_int2;
  assign restfa2_in13_int0 = restfa_in10_c ^ restfa_in11_c;
  assign restfa2_in13_int1 = restfa_in10_c & restfa_in11_c;
  assign restfa2_in13_int2 = restfa1_in13_c & restfa2_in13_int0;
  assign restfa2_in13_s = restfa2_in13_int0 ^ restfa1_in13_c;
  assign restfa2_in13_c = restfa2_in13_int1 | restfa2_in13_int2;
  
  
  
   
  
  assign rest_in14_s = rest_in12_s ^ rest_in13_s;
  assign rest_in14_c = rest_in12_s & rest_in13_s;
  assign restfa1_in14_int0 = restfa1_in12_s ^ restfa1_in13_s;
  assign restfa1_in14_int1 = restfa1_in12_s & restfa1_in13_s;
  assign restfa1_in14_int2 = rest_in14_c & restfa1_in14_int0;
  assign restfa1_in14_s = restfa1_in14_int0 ^ rest_in14_c;
  assign restfa1_in14_c = restfa1_in14_int1 | restfa1_in14_int2;
  assign restfa2_in14_int0 = restfa2_in12_s ^ restfa2_in13_s;
  assign restfa2_in14_int1 = restfa2_in12_s & restfa2_in13_s;
  assign restfa2_in14_int2 = restfa1_in14_c & restfa2_in14_int0;
  assign restfa2_in14_s = restfa2_in14_int0 ^ restfa1_in14_c;
  assign restfa2_in14_c = restfa2_in14_int1 | restfa2_in14_int2;
  assign restfa3_in14_int0 = restfa2_in12_c ^ restfa2_in13_c;
  assign restfa3_in14_int1 = restfa2_in12_c & restfa2_in13_c;
  assign restfa3_in14_int2 = restfa2_in14_c & restfa3_in14_int0;
  assign restfa3_in14_s = restfa3_in14_int0 ^ restfa2_in14_c;
  assign restfa3_in14_c = restfa3_in14_int1 | restfa3_in14_int2;





  assign rest = (~restfa3_in14_c) & (~restfa3_in14_s) & (~restfa2_in14_s) & (~restfa1_in14_s) & rest_in14_s;
  //assign rest = (~restfa3_in14_c) & (~restfa3_in14_s) & (~restfa2_in14_s) & (restfa1_in14_s) & (~rest_in14_s);
  //assign rest = (~restfa3_in14_c) & (~restfa3_in14_s) & (~restfa2_in14_s) & (restfa1_in14_s) & rest_in14_s;



  assign po11 = po11_prelocked ^ hd ^ rest;
  assign po12 = po12_prelocked ^ hd ^ rest;
  assign po13 = po13_prelocked ^ hd ^ rest;
  assign po14 = po14_prelocked ^ hd ^ rest;
  assign po15 = po15_prelocked ^ hd ^ rest;
  assign po16 = po16_prelocked ^ hd ^ rest;
  assign po17 = po17_prelocked ^ hd ^ rest;
  assign po18 = po18_prelocked ^ hd ^ rest;
  assign po19 = po19_prelocked ^ hd ^ rest;
  assign po20 = po20_prelocked ^ hd ^ rest;
  assign po21 = po21_prelocked ^ hd ^ rest;

endmodule


